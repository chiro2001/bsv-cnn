import FixedPoint::*;

typedef 28 InputHeight;
typedef 28 InputWidth;
typedef FixedPoint#(12, 20) ElementType;