import Data::*;

module mkTb();

endmodule