import FixedPoint::*;

typedef 28 InputHeight;
typedef 28 InputWidth;
// 32bits
// typedef FixedPoint#(12, 20) ElementType;
// 16bits
typedef FixedPoint#(6, 10) ElementType;

typedef Bit#(4) ResultType;