import FIFOF::*;
import Vector::*;
import Data::*;

interface Layer#(type in, type out);
  method Action put(in x);
  method ActionValue#(out) get;
endinterface

module mkFCLayer#(parameter String layer_name)(Layer#(in, out))
  provisos(
    Bits#(out, lines_bits), 
    Bits#(in, depth_bits), 
    Mul#(lines, 8, lines_bits), 
    Mul#(depth, 8, depth_bits),
    PrimSelectable#(in, Int#(8)),
    PrimSelectable#(out, Int#(8)),
    PrimWriteable#(Reg#(out), Int#(8))
  );
  LayerData_ifc#(Int#(8), lines, depth) data <- mkLayerData(layer_name);
  Reg#(Bool) stage <- mkReg(False);
  Reg#(Bool) done <- mkReg(True);
  Reg#(out) tmp <- mkReg(unpack('0));

  FIFOF#(in) fifo_in <- mkFIFOF1;
  FIFOF#(out) fifo_out <- mkFIFOF1;

  rule start (!stage && done && data.weightsDone() && data.biasDone());
    $display("Layer %s start", layer_name);
    data.weightStart();
    done <= False;
    tmp <= unpack('0);
  endrule

  rule acc_weights (!stage && !done && !data.weightsDone() && data.biasDone());
    let index = data.getIndex() - 1;
    // $display("Layer %s acc weights, index=%x", layer_name, index);
    let weight = data.getWeight();
    let top = fifo_in.first;
    out t = tmp;
    for (Integer i = 0; i < valueOf(lines); i = i + 1) begin
      let w <- weight[i];
      let mul = top[i] * w;
      t[i] = tmp[i] + (mul >> 6);
    end
    tmp <= t;
  endrule

  rule acc_weights_to_bias (!stage && !done && data.weightsDone() && data.biasDone());
    // $display("Layer %s acc weights to bias", layer_name);
    data.biasStart();
    stage <= True;
  endrule

  rule acc_bias (stage && !done && data.weightsDone() && !data.biasDone());
    let index_bias = data.getIndexLines() - 1;
    // $display("Layer %s acc bias, index_bias=%x", layer_name, index_bias);
    let bias <- data.getBias();
    out t = tmp;
    t[index_bias] = tmp[index_bias] + bias;
    tmp <= t;
  endrule

  rule acc_bias_to_fifo_out (stage && !done && data.weightsDone() && data.biasDone());
    // $display("Layer %s acc bias to fifo out", layer_name);
    done <= True;
  endrule

  rule do_fifo_out (stage && done && data.weightsDone() && data.biasDone());
    // $display("Layer %s do fifo out", layer_name);
    fifo_out.enq(tmp);
    fifo_in.deq;
    stage <= False;
    tmp <= unpack('0);
  endrule

  method Action put(in x);
    fifo_in.enq(x);
  endmethod

  method ActionValue#(out) get;
    out y = fifo_out.first;
    fifo_out.deq;
    return y;
  endmethod
endmodule