// import Float32::*;

module mkTb();

  // FpPairIfc#(32) mult <- mkFpMult32;

  rule test_mult;
    $display("no floating point support yet");
    $finish;
  endrule
endmodule
