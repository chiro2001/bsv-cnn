import Float32::*;

module mkTb();

endmodule