// import Float32::*;

module mkTb();

  // FpPairIfc#(32) mult <- mkFpMult32;

  rule test_mult;
    
  endrule
endmodule
